moudule 
begin
end
endmodule
