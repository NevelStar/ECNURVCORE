
module edge_detector
(
	input		rst_n,
	input		clk,
	input		level_i,
	output		edge_o
	
);